   ������2D:\DSNetworkS\DSN_Structure\usr\bin\pRaport8v3.exe����� ������:D:\DSNetworkS\DSN_Structure\usr\bin\pOreolVolumeReset3.exe��������� �������5D:\DSNetworkS\DSN_Structure\usr\bin\pOreolSetTime.exeNoItem 3NoPath 3NoItem 4NoPath 4NoItem 5NoPath 5NoItem 6NoPath 6NoItem 7NoPath 7NoItem 8NoPath 8NoItem 9NoPath 9                pB   A  P4Db@  P`(�?              pB   A  P4Db@  P`(�?              pB   A  P4Db@  P`(�?              pB   A  P4Db@  P`(�?              pB   A  P4Db@  P`(�?   :                         d       