      $@      4@      Y@      @      $@      Y@����              >@      >@      0@                     �r@      @      Y@      4@     �A@   ����?   ����?   �̬Q@                      �?      $@                              �?    �����	�������������1�������2D:\DSNetwork\DSN_Structure\usr\bin\KBI20090605.xls                                                                         ��@                 ������.\pRaport9.exe����� �� ��.\pOreolSetTime.exe����� ������.\pOreolVolumeReset.exe
����������.\pOreolSetBlock.exe����� ���������.\pOreolRestart.exepOreolVolumeReset3#E:\Oreol\bin\pOreolVolumeReset3.exeNoItem 6NoPath 6NoItem 7NoPath 7NoItem 8NoPath 8NoItem 9NoPath 9                  ��F   A  0�)�?  (h0� @              pB   A  ��tf@  (h0� @              �D   A  `�'�@  (h0� @              �C   A  `�'�=@  (h0� @              �D   A  �>G"@  (h0� @   �   �  