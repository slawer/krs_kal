      $@      4@      Y@      @      $@      Y@����              >@      >@      0@                     �r@      @      Y@      4@     �A@   ����?   ����?   �̬Q@                      �?      $@                              �?    �����������2���12D:\DSNetwork\DSN_Structure\usr\bin\KBI20090605.xls                                                                                               NoItem 0NoPath 0NoItem 1NoPath 1NoItem 2NoPath 2NoItem 3NoPath 3NoItem 4NoPath 4NoItem 5NoPath 5NoItem 6NoPath 6NoItem 7NoPath 7NoItem 8NoPath 8NoItem 9NoPath 9                  4E   A  �@  (h0� @              pC   A  P4DB@  (h0� @             ��F   A  Ѓ�H�?  (h0� @              �B   A  P4DR@  (h0� @               4E   A   @铦?  (h0� @   �   �  