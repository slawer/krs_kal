      $@      4@      Y@      @      $@      Y@����              >@      >@      .@      @      @     �r@      @      Y@      4@     �K@   ����?   ����?  �,3�l@                      I@      I@                             �?    ����������������_����������������
C:\KBI.xls                                                                                              ����� ������:D:\DSNetworkS\DSN_Structure\usr\bin\pOreolVolumeReset3.exe��������� �������5D:\DSNetworkS\DSN_Structure\usr\bin\pOreolSetTime.exeRaport9>D:\DSNetworkS\DSN_Structure\usr\bin\pRaport9v2_101102_1742.exefilter.D:\DSNetworkS\DSN_Structure\usr\bin\filter.exepOreolVolumeReset3#D:\Oreol\bin\pOreolVolumeReset3.exepOreolSetBlockD:\Oreol\bin\pOreolSetBlock.exepOreolSetTime2D:\Oreol\bin\pOreolSetTime2.exe�������D:\Oreol\bin\pOreolRestart.exeNoItem 8NoPath 8NoItem 9NoPath 9                  4E   A  �>G@  <*��?                pB   A  ���jk@   ඬ�?              �D   A  �bd-@   ඬ�?               4D   A  �bd=@  <*��?               4E   A  `�'�@  <*��?   �   %  