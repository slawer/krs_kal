      $@      4@      Y@      @      $@      Y@����              >@      >@      0@                     �r@      @      Y@      4@     �A@   ����?   ����?   �̬Q@                      �?      $@                              �?    �����614-2168��351722D:\DSNetwork\DSN_Structure\usr\bin\KBI20090605.xls                                                                        ��@                 ����� ������#C:\Oreol\bin\pOreolVolumeReset3.exe����C:\Oreol\bin\pOreolSetTime.exepRaport9C:\Oreol\bin\pRaport9.exeNoItem 3NoPath 3NoItem 4NoPath 4NoItem 5NoPath 5NoItem 6NoPath 6NoItem 7NoPath 7NoItem 8NoPath 8NoItem 9NoPath 9                   �B   A  ���b@  (h0� @                 �B   A  ���c@  (h0� @                 4D   A  ��7@  (h0� @                 �C   A  ��G@  (h0� @                 pB   A  �L�q@  (h0� @    �   %  